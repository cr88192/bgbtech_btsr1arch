/*
Detect unconditional branch instructions for early branch.
Happens in parallel with the main ID1 stage.

May also incorporate branch prediction.

exBraDir:
* (1:0) = Branch Direction (Predication Mode)
** 00: Unconditional
** 01: Not a Branch
** 10: Branch if True
** 11: Branch if False
* (  2) = Branch was not taken

State of Branch:
* 000: Branch not taken (Weak)
* 011: Branch not taken (Strong)
* 100: Branch taken (Strong)
* 111: Branch taken (Weak)

State Machine 2:
* 000: Weak Not Taken			(0->001, 1->110)
* 001: Strong Not Taken			(0->001, 1->000)
* 010: Trans Weak, Not Taken	(0->000, 1->111)
* 011: Trans Strong, Not Taken	(0->010, 1->111)
* 100: Weak Taken				(0->010, 1->101)
* 101: Strong Taken				(0->100, 1->101)
* 110: Trans Weak, Taken		(0->011, 1->100)
* 111: Trans Strong, Taken		(0->011, 1->110)

*/

module DecPreBra(
	clock,		reset,
	istrWord,	istrBasePc,	istrBraPc,
	preBraPc,	preIsBra,
	regValLr,	ifBraBPc,
	exBraBPc,	exBraDir);

input			clock;
input			reset;
input[63:0]		istrWord;	//Instruction Word
input[47:0]		istrBasePc;	//Instruction Base PC
input[47:0]		istrBraPc;	//Branch Base PC
input[63:0]		regValLr;	//Link Register

input[47:0]		ifBraBPc;	//Fetch Branch PC
input[47:0]		exBraBPc;	//Fetch Base PC
input[2:0]		exBraDir;

output[47:0]	preBraPc;
output			preIsBra;

reg[47:0]	tPreBraPc;
reg			tPreBra;
assign	preBraPc	= tPreBraPc;
assign	preIsBra	= tPreBra;


// reg[32:0]	tBraDisp8;
// reg[32:0]	tBraDisp20;
reg[24:0]	tBraDisp8;
reg[24:0]	tBraDisp20;

reg[31:0]	tDisp8;
reg[31:0]	tDisp20;

reg[11:0]	tBraDisp8HiP0;
reg[11:0]	tBraDisp8HiP1;
reg[11:0]	tBraDisp8HiN1;

reg[20:0]	tBraDisp8Lo;
reg[20:0]	tBraDisp20Lo;

reg			tIsBra8;		//Unconditional Branch (8-bit Disp)
reg			tIsBra20;		//Unconditional Branch (16-bit Disp)
reg			tIsRtsu;

reg			tIsBraCc8;		//Conditional Branch (8-bit Disp)
reg			tIsBraCc20;		//Conditional Branch (20-bit Disp)
reg			tDoBraCc8;		//Take Conditional Branch (Cc8)
reg			tDoBraCc20;		//Take Conditional Branch (Cc20)

reg[2:0]	preCnts[63:0];
// reg[2:0]	preCnts[4095:0];
reg[2:0]	tPreIfCnt;
reg[2:0]	tPreExCnt;
reg[2:0]	tPreExCntB;
reg[2:0]	tPreExDir;
reg[47:0]	tPreExBPc;

// reg[5:0]	preBits[63:0];
reg[5:0]	tPreIfBit;
reg[5:0]	tPreExBit;
reg[5:0]	tPreExBitB;
reg			tPreBit;

reg[5:0]	tPreIfIx;
reg[5:0]	tPreIdIx;
reg[5:0]	tPreIbIx;
reg[5:0]	tPreExIx;
reg[5:0]	tPreExIxA;

//reg[11:0]	tPreIfIx;
//reg[11:0]	tPreIdIx;
//reg[11:0]	tPreIbIx;
//reg[11:0]	tPreExIx;
//reg[11:0]	tPreExIxA;

reg[5:0]	tHistBits;
reg[5:0]	tHistBitsB;

always @*
begin
//	tPreBraPc	= UV48_XX;
	tPreBraPc	= istrBraPc;
	tPreBra		= 0;
	tHistBitsB	= tHistBits;
	
	tPreIfIx	= ifBraBPc[6:1]		^ tHistBits;
	tPreIbIx	= istrBasePc[6:1]	^ tHistBits;
	tPreExIxA	= exBraBPc[6:1]		^ tHistBits;

//	tPreIfIx	= ifBraBPc[12:1];
//	tPreIbIx	= istrBasePc[12:1];
//	tPreExIxA	= exBraBPc[12:1];
	
	tPreExCntB	= tPreExCnt;
	tPreExBitB	= tPreExBit;

	if(tPreExDir[1])
	begin
		tHistBitsB = { tHistBits[4:0], tPreExDir[2] };
		tPreExBitB = { tPreExBit[4:0], tPreExDir[2] };

		case( {tPreExDir[2], tPreExCnt[2:0]} )
			4'b0000: tPreExCntB=3'b001;
			4'b0001: tPreExCntB=3'b001;
			4'b0010: tPreExCntB=3'b000;
			4'b0011: tPreExCntB=3'b010;
			4'b0100: tPreExCntB=3'b010;
			4'b0101: tPreExCntB=3'b100;
			4'b0110: tPreExCntB=3'b011;
			4'b0111: tPreExCntB=3'b011;
			4'b1000: tPreExCntB=3'b110;
			4'b1001: tPreExCntB=3'b000;
			4'b1010: tPreExCntB=3'b111;
			4'b1011: tPreExCntB=3'b111;
			4'b1100: tPreExCntB=3'b101;
			4'b1101: tPreExCntB=3'b101;
			4'b1110: tPreExCntB=3'b100;
			4'b1111: tPreExCntB=3'b110;
		endcase

//		$display("PreBra: Predict State %X, BPc=%X",
//			{tPreExDir[2], tPreExCnt[2:0]},
//			tPreExBPc);
	end
		
	tDisp8		= { istrWord[7]?UV24_FF:UV24_00, istrWord[7:0] };
	tDisp20		= {
		istrWord[7]?UV12_FF:UV12_00,
		istrWord[7:0], istrWord[27:16] };
	
//	tBraDisp8	= {1'b0, istrBraPc[31:0] } + { tDisp8[31:0], 1'b0 };
//	tBraDisp20	= {1'b0, istrBraPc[31:0] } + { tDisp20[31:0], 1'b0 };
	tBraDisp8	= {1'b0, istrBraPc[23:0] } + { tDisp8[23:0], 1'b0 };
	tBraDisp20	= {1'b0, istrBraPc[23:0] } + { tDisp20[23:0], 1'b0 };

// `ifdef def_true
`ifndef def_true
	tBraDisp8HiP0	= istrBraPc[31:21];
	tBraDisp8HiP1	= istrBraPc[31:21]+1;
	tBraDisp8HiN1	= istrBraPc[31:21]-1;
	tBraDisp8Lo		= { 1'b0, istrBraPc[20:1]} + tDisp8[19:0];
	tBraDisp20Lo	= { 1'b0, istrBraPc[20:1]} + tDisp20[19:0];

	if(tDisp8[30])
		tBraDisp8 = {
			tBraDisp8Lo[20] ? tBraDisp8HiP0 : tBraDisp8HiN1,
			tBraDisp8Lo[19:0], istrBraPc[0]	};
	else
		tBraDisp8 = {
			tBraDisp8Lo[20] ? tBraDisp8HiP1 : tBraDisp8HiP0,
			tBraDisp8Lo[19:0], istrBraPc[0]	};

	if(tDisp20[30])
		tBraDisp20 = {
			tBraDisp20Lo[20] ? tBraDisp8HiP0 : tBraDisp8HiN1,
			tBraDisp20Lo[19:0], istrBraPc[0]	};
	else
		tBraDisp20 = {
			tBraDisp20Lo[20] ? tBraDisp8HiP1 : tBraDisp8HiP0,
			tBraDisp20Lo[19:0], istrBraPc[0]	};
`endif

	tIsBra8		=
		(istrWord[15:12]==4'h2) &&
		(istrWord[11: 9]==3'b000);
//		(istrWord[11: 8]==4'b0000);
	tIsBra20		=
		(istrWord[15:12]==4'hF) &&
		(istrWord[11: 8]==4'h0) &&
		(istrWord[31:29]==3'b110);
//		(istrWord[31:28]==4'b1100);

	tIsBraCc8		=
		(istrWord[15:12]==4'h2) &&
		(istrWord[11: 9]==3'b001);
	tIsBraCc20		=
		(istrWord[15:12]==4'hF) &&
		(istrWord[11: 8]==4'h0) &&
		(istrWord[31:29]==3'b111);
	
	tIsRtsu			=
		(istrWord[15:0] == 16'h3012);

//	tIsBra8		= 0;
//	tIsBra20	= 0;
//	tIsRtsu		= 0;

	tDoBraCc8	= 0;
	tDoBraCc20	= 0;

// `ifndef def_true
`ifdef def_true
	if(tIsBraCc8 && (tPreIbIx==tPreIdIx))
	begin
//		tDoBraCc8 = tPreExCntB[1] ? tPreBit : tPreIfCnt[2];
		tDoBraCc8 = tPreIfCnt[2] ^ tPreIfCnt[1];
		
//		tDoBraCc8 = tPreBit;
//		tDoBraCc8 = tPreIfCnt[2];
//		tDoBraCc8 = !tPreIfCnt[2];
//		$display("PreBra: Predict 8, Do=%d, BPc=%X",
//			tDoBraCc8, istrBasePc);
	end

	if(tIsBraCc20 && (tPreIbIx==tPreIdIx))
	begin
//		tDoBraCc20 = tPreExCntB[1] ? tPreBit : tPreIfCnt[2];
		tDoBraCc20 = tPreIfCnt[2] ^ tPreIfCnt[1];
		
//		tDoBraCc20 = tPreBit;
//		tDoBraCc20 = tPreIfCnt[2];
//		tDoBraCc20 = !tPreIfCnt[2];
//		$display("PreBra: Predict 20, Do=%d", tDoBraCc20);
	end
`endif
	
	if(tIsBra8 || tIsBraCc8)
	begin
//		tPreBraPc	= { istrBraPc[47:32], tBraDisp8[31:0] };
		tPreBraPc	= { istrBraPc[47:24], tBraDisp8[23:0] };
	end

	if(tIsBra20 || tIsBraCc20)
	begin
//		tPreBraPc	= { istrBraPc[47:32], tBraDisp20[31:0] };
		tPreBraPc	= { istrBraPc[47:24], tBraDisp20[23:0] };
	end

//	if(tIsBra8)
	if(tIsBra8 || tDoBraCc8)
	begin
//		$display("PreBra: BRA8, PC=%X I=%X-%X PC2=%X",
//			istrBasePc,
//			istrWord[15:0], istrWord[31:16],
//			tBraDisp8);
//		tPreBraPc	= tBraDisp8;
//		tPreBraPc	= { istrBraPc[47:32], tBraDisp8 };
		tPreBra		= 1;
		
//		if(tBraDisp8[32])
		if(tBraDisp8[24])
			tPreBra		= 0;
	end

//	if(tIsBra20)
	if(tIsBra20 || tDoBraCc20)
	begin
//		$display("PreBra: BRA20, I=%X-%X PC2=%X",
//			istrWord[15:0], istrWord[31:16], tBraDisp20);
//		tPreBraPc	= tBraDisp20;
//		tPreBraPc	= { istrBraPc[47:32], tBraDisp20 };
		tPreBra		= 1;

//		if(tBraDisp20[32])
		if(tBraDisp20[24])
			tPreBra		= 0;
	end
	
	if(tIsRtsu)
	begin
//		$display("PreBra: RTSU, I=%X-%X PC2=%X",
//			istrWord[15:0], istrWord[31:16], regValLr);
		tPreBraPc	= regValLr[47:0];
		tPreBra		= 1;
	end

//	tPreBra		= 0;
end

always @(posedge clock)
begin
	tHistBits	<= tHistBitsB;
	tPreExBit	<= tPreExBitB;

	tPreIfCnt	<= preCnts[tPreIfIx];
	tPreIdIx	<= tPreIfIx;

	tPreExCnt			<= preCnts[tPreExIxA];
	preCnts[tPreExIx]	<= tPreExCntB;
	tPreExIx			<= tPreExIxA;
	tPreExDir			<= exBraDir;
	tPreExBPc			<= exBraBPc;
end

endmodule